library verilog;
use verilog.vl_types.all;
entity test_send_sv_unit is
end test_send_sv_unit;
