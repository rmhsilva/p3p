library verilog;
use verilog.vl_types.all;
entity test_gdp_controller_sv_unit is
end test_gdp_controller_sv_unit;
