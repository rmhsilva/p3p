library verilog;
use verilog.vl_types.all;
entity top_level_sv_unit is
end top_level_sv_unit;
