library verilog;
use verilog.vl_types.all;
entity max_sv_unit is
end max_sv_unit;
