library verilog;
use verilog.vl_types.all;
entity test_top_level_sv_unit is
end test_top_level_sv_unit;
