library verilog;
use verilog.vl_types.all;
entity test_gdp is
end test_gdp;
