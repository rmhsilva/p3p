library verilog;
use verilog.vl_types.all;
entity test_send is
end test_send;
