library verilog;
use verilog.vl_types.all;
entity send_sv_unit is
end send_sv_unit;
