library verilog;
use verilog.vl_types.all;
entity all_s_data_sv_unit is
end all_s_data_sv_unit;
