library verilog;
use verilog.vl_types.all;
entity sram_sv_unit is
end sram_sv_unit;
