library verilog;
use verilog.vl_types.all;
entity gdp_controller_sv_unit is
end gdp_controller_sv_unit;
