library verilog;
use verilog.vl_types.all;
entity test_top_level is
end test_top_level;
