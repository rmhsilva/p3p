library verilog;
use verilog.vl_types.all;
entity test_uart_sv_unit is
end test_uart_sv_unit;
