library verilog;
use verilog.vl_types.all;
entity test_uart is
end test_uart;
