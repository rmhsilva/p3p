library verilog;
use verilog.vl_types.all;
entity gdp_sv_unit is
end gdp_sv_unit;
