library verilog;
use verilog.vl_types.all;
entity uart_sv_unit is
end uart_sv_unit;
