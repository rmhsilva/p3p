library verilog;
use verilog.vl_types.all;
entity normaliser_sv_unit is
end normaliser_sv_unit;
